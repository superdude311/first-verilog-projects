// testbench for 6502 multiplication accelerator

module tb;
    timeunit 1ns;
    timeprecision 1ps;

    logic clk;
    logic RWB;
    logic CE;
    logic A0;
    logic [7:0] A;
    logic [7:0] B;
    logic [7:0] Dout;
    logic [15:0] out;
    wire [7:0] D;
    



endmodule